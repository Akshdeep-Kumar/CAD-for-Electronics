** Profile: "SCHEMATIC1-DC_analysis"  [ C:\Users\akshd\Documents\MAIN\Extras\CAD_Lab_self\E1-PSpiceFiles\SCHEMATIC1\DC_analysis.sim ] 

** Creating circuit file "DC_analysis.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\akshd\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0v 5v 0.1v 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
